`timescale 1ns / 1ps

////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer:
//
// Create Date:   14:22:15 01/31/2014
// Design Name:   writeback
// Module Name:   /home/pravinkumar/Workspace/Xilinx/AsynARM/writeback_test.v
// Project Name:  arm
// Target Device:  
// Tool versions:  
// Description: 
//
// Verilog Test Fixture created by ISE for module: writeback
//
// Dependencies:
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
////////////////////////////////////////////////////////////////////////////////

module writeback_test;
//
//	// Outputs
//	wire ;
//
//	// Instantiate the Unit Under Test (UUT)
//	writeback uut (
//		.()
//	);
//
//	initial begin
//		// Initialize Inputs
//
//		// Wait 100 ns for global reset to finish
//		#100;
//        
//		// Add stimulus here
//
//	end
      
endmodule

